`define B115200 868
`define B57600 1736
`define B38400 2604
`define B19200 5208
`define B9600 10417
`define B4800 20833
`define B2400 41667
`define B1200 83333
`define B600 166667
`define B300 333333
