// Top module

module blank (
  input clk_100mhz
);

endmodule
